module fir_handle
(
	output sink_valid,
	output sink_ready
);

assign sink_valid=1'b1;
assign sink_ready=1'b1;

endmodule 